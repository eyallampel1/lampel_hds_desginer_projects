--
-- VHDL Architecture my_project_lib.HexTimer.behave
--
-- Created:
--          by - Suzana.UNKNOWN (SUZANA-PC)
--          at - 21:15:04 27/02/2016
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY HexTimer IS
   PORT( 
      clk25          : IN     std_logic;
      somePushButton : IN     std_logic
   );

-- Declarations

END HexTimer ;

--
ARCHITECTURE behave OF HexTimer IS
BEGIN
END behave;

